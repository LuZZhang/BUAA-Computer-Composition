`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   10:18:31 12/14/2017
// Design Name:   mips
// Module Name:   D:/jizu/homework/P4_plus/P4_plus/tb.v
// Project Name:  P4_plus
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: mips
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module tb;

	// Inputs
	reg clk;
	reg reset;

	// Instantiate the Unit Under Test (UUT)
	mips uut (
		.clk(clk), 
		.reset(reset)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 1;
		# 10;
      reset = 0;
		// Wait 100 ns for global reset to finish
		
        
		// Add stimulus here

	end
      always #5 clk = ~clk;
endmodule

